//  Module: and_module.sv
//qualcosa li

module and_module.sv
    (
        input logic a,
        input logic b,
        output logic y
    );

    assign y = a + b;
endmodule: and_module.sv
